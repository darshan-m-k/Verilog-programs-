module multiplier_tb();
  reg [3:0]a;
  wire [6:0]y1,y2;
  multi8 dut(a,y1,y2);
  initial begin
    a=4'b0000;  #10
    a=4'b0010;  #10
    a=4'b0100;  #10
    a=4'b0110;  #10;
  end
  initial begin 
    $monitor ( " sim time = %t, a=%b, 
y1=%b, y2=%b", $time,a,y1,y2);
  end
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0,a,y1,y2);
  end 
endmodule

*************************************DESIGN CODE*****************************

// Dataflow Modelling

module majority_1(A,B,C,F);
  input A,B,C;
  output F;
  assign F = (A&B)|(A&C)|(B&C);
endmodule

//Gatelevel Modelling

module majority_1(A,B,C,F);
  input A,B,C;
  output F;
  wire w1,w2,w3;
  and a1(w1,B,C);
  and a2(w2,A,C);
  and a3(w3,A,B);
  or o1(F,w1,w2,w3);
endmodule

/////////////////////////////////////////////////////////////////

***********************************TESTBENCH*************************************

module tb_majority_1;
  reg A, B, C;
  wire F;
  majority_1 DUT(A,B,C,F);
  initial begin
        A = 1'b0; B = 1'b0; C = 1'b0; 
    #10;    A = 1'b0; B = 1'b0; C = 1'b1;
    #10;    A = 1'b0; B = 1'b1; C = 1'b0; 
    #10; 	A = 1'b0; B = 1'b1; C = 1'b1;
    #10;    A = 1'b1; B = 1'b0; C = 1'b0;
    #10;    A = 1'b1; B = 1'b0; C = 1'b1; 
    #10;    A = 1'b1; B = 1'b1; C = 1'b0;
    #10;    A = 1'b1; B = 1'b1; C = 1'b1;
  end
  initial begin 
   $monitor("simtime=%0t,A=%b,B=%b,C=%b,F=%b",$time,A,B,C,F);
  end
	initial begin 
     $dumpfile("dump.vcd");
     $dumpvars(0,A,B,C,F);
    end  
endmodule
